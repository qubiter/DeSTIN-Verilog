`timescale 1ns / 100ps

module starveunit()
  
endmodule